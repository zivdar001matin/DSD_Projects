ENTITy alu_tb IS
END alu_tb;
