
-- g_<name> corresponds to Generic
-- p_<name> corresponds to Port
-- c_<name> corresponds to Constant
-- s_<name> corresponds to Signal

-- Packages
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

-- Entity Port and Generic
ENTITY alu IS 
    GENERIC (
        g_size : integer := 32
    );
    PORT(
        p_A     : IN signed(g_size - 1 DOWNTO 0);
        p_B     : IN signed(g_size - 1 DOWNTO 0);
        p_cin   : IN integer;
        p_sin   : IN std_logic;
        p_funct : IN signed(3 DOWNTO 0);
        p_sout  : OUT std_logic;
        p_cout  : OUT std_logic;
        p_Ov    : OUT std_logic;
        p_Z     : OUT signed(g_size - 1 DOWNTO 0)
    );
END alu;

-- Entity Architecture
ARCHITECTURE arch OF alu IS
    -- Design decision
    CONSTANT c_zero : signed(g_size -1 DOWNTO 0) := (others => '0');

    SIGNAL s_AplusB         : signed(g_size DOWNTO 0);
    SIGNAL s_AplusBplusCin  : signed(g_size DOWNTO 0);

BEGIN
    s_AplusB <= ('0' & p_A) + ('0' & p_B);
    s_AplusBplusCin <= ('0' & p_A) + ('0' & p_B) + p_cin;
    PROCESS(p_A, p_B, p_cin, p_sin, p_funct)
    BEGIN
        IF p_funct = "0000" THEN
            p_Z <= NOT p_B(g_size - 1) & p_B(g_size - 2 DOWNTO 0);
        ELSIF p_funct = "0001" THEN
            p_Z <= s_AplusB(g_size - 1 DOWNTO 0);
            p_cout <= s_AplusB(g_size);
            p_Ov <= (p_A(g_size - 1) AND p_B(g_size - 1) AND NOT s_AplusB(g_size - 1)) OR
                (NOT p_A(g_size - 1) AND NOT p_B(g_size - 1) AND s_AplusB(g_size - 1));
        ELSIF p_funct = "0010" THEN
            p_Z <= s_AplusBplusCin(g_size - 1 DOWNTO 0);
            p_cout <= s_AplusBplusCin(g_size);
            p_Ov <= (p_A(g_size - 1) AND p_B(g_size - 1) AND NOT s_AplusBplusCin(g_size - 1)) OR
                (NOT p_A(g_size - 1) AND NOT p_B(g_size - 1) AND s_AplusBplusCin(g_size - 1));
        ELSIF p_funct = "0011" THEN
            p_Z <= p_A - p_B;
        ELSIF p_funct = "0100" THEN
            p_Z <= -p_B;
        ELSIF p_funct = "0101" THEN
            p_Z <= NOT p_B;
        ELSIF p_funct = "0110" THEN
            p_Z <= p_A AND p_B;
        ELSIF p_funct = "0111" THEN
            p_Z <= p_A OR p_B;
        ELSIF p_funct = "1000" THEN
            p_Z <= p_A XOR p_B;
        ELSIF p_funct = "1001" THEN
            p_Z <= p_A(g_size  - 2 DOWNTO 0) & p_sin;
            p_sout <= p_A(g_size  - 1);
        ELSIF p_funct = "1010" THEN
            p_Z <= p_sin & p_A(g_size  - 1 DOWNTO 1);
            p_sout <= p_A(0);
        ELSIF p_funct = "1011" THEN
            p_Z <= p_A rol 1;
        ELSIF p_funct = "1100" THEN
            p_Z <= p_A ror 1;
        ELSIF p_funct = "1101" THEN
            IF p_A > p_B THEN
                p_Z <= c_zero + 1;
            ELSE
                p_Z <=  c_zero;
            END IF;
        ELSIF p_funct = "1110" THEN
            IF p_A < p_B THEN
                p_Z <= c_zero + 1;
            ELSE
                p_Z <= c_zero;
            END IF;
        ELSIF p_funct = "1111" THEN
            IF p_A = p_B THEN
                p_Z <= c_zero + 1;
            ELSE
                p_Z <= c_zero;
            END IF;
        ELSE
            p_Z <= c_zero;
        END IF;
    END PROCESS;
END arch;